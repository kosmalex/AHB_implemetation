package util;
  typedef enum logic[1:0] {IDLE, BUSY, NONSEQ, SEQ} trans_t;
endpackage